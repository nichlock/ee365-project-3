-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version
-- Created on Tue Oct 12 16:30:18 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY encoder_sm IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        a : IN STD_LOGIC := '0';
        b : IN STD_LOGIC := '0';
        add : OUT STD_LOGIC;
        sub : OUT STD_LOGIC
    );
END encoder_sm;

ARCHITECTURE BEHAVIOR OF encoder_sm IS
    TYPE type_fstate IS (init,from_left,from_right,in_middle_from_left,in_middle_from_right,leaving_from_left,leaving_from_right,add_one,sub_one);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,a,b)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= init;
            add <= '0';
            sub <= '0';
        ELSE
            add <= '0';
            sub <= '0';
            CASE fstate IS
                WHEN init =>
                    IF (((a = '1') AND NOT((b = '1')))) THEN
                        reg_fstate <= from_left;
                    ELSIF ((NOT((a = '1')) AND (b = '1'))) THEN
                        reg_fstate <= from_right;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= init;
                    END IF;
                WHEN from_left =>
                    IF (((a = '1') AND (b = '1'))) THEN
                        reg_fstate <= in_middle_from_left;
                    ELSIF (((a = '1') AND NOT((b = '1')))) THEN
                        reg_fstate <= from_left;
                    ELSE
                        reg_fstate <= init;
                    END IF;
                WHEN from_right =>
                    IF (((a = '1') AND (b = '1'))) THEN
                        reg_fstate <= in_middle_from_right;
                    ELSIF (((b = '1') AND NOT((a = '1')))) THEN
                        reg_fstate <= from_right;
                    ELSE
                        reg_fstate <= init;
                    END IF;
                WHEN in_middle_from_left =>
                    IF ((NOT((a = '1')) AND (b = '1'))) THEN
                        reg_fstate <= leaving_from_left;
                    ELSIF (((a = '1') AND (b = '1'))) THEN
                        reg_fstate <= in_middle_from_left;
                    ELSE
                        reg_fstate <= init;
                    END IF;
                WHEN in_middle_from_right =>
                    IF (((a = '1') AND NOT((b = '1')))) THEN
                        reg_fstate <= leaving_from_right;
                    ELSIF (((a = '1') AND (b = '1'))) THEN
                        reg_fstate <= in_middle_from_right;
                    ELSE
                        reg_fstate <= init;
                    END IF;
                WHEN leaving_from_left =>
                    IF ((NOT((a = '1')) AND NOT((b = '1')))) THEN
                        reg_fstate <= add_one;
                    ELSIF ((NOT((a = '1')) AND (b = '1'))) THEN
                        reg_fstate <= leaving_from_left;
                    ELSE
                        reg_fstate <= init;
                    END IF;
                WHEN leaving_from_right =>
                    IF ((NOT((a = '1')) AND NOT((b = '1')))) THEN
                        reg_fstate <= sub_one;
                    ELSIF ((NOT((b = '1')) AND (a = '1'))) THEN
                        reg_fstate <= leaving_from_right;
                    ELSE
                        reg_fstate <= init;
                    END IF;
                WHEN add_one =>
                    reg_fstate <= init;

                    add <= '1';
                WHEN sub_one =>
                    reg_fstate <= init;

                    sub <= '1';
                WHEN OTHERS => 
                    add <= 'X';
                    sub <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
